/**
 * name: alu.sv
 * desc: 
 */

module ALU (
    input   logic [3:0]     ctrl,
    input   logic [31:0]    arg1,
    input   logic [31:0]    arg2,
    output  logic           zero        = 'd0, // zero or not
    output  logic [31:0]    result      = 32'd0 
);
    /* ctrls */
    parameter ctrl_addiu    = 4'b0000;
    parameter ctrl_sw       = 4'b0001;
    parameter ctrl_addu     = 4'b0010;
    parameter ctrl_invalid  = 4'bxxxx;

    always_comb 
        case (ctrl)
            /* addiu */
            ctrl_addiu: begin
                zero    = arg1 == arg2 ? 1'b1 : 1'b0;
                result  = arg1 + arg2;
            end
            /* sw */
            ctrl_sw: begin
                zero    = arg1 == arg2 ? 1'b1 : 1'b0;
                result  = arg1 + arg2;
            end
            /* addu */
            ctrl_addu: begin
                zero    = arg1 == arg2 ? 1'b1 : 1'b0;
                result  = arg1 + arg2;
            end
            default: begin
                zero    = 1'bx;
                result  = 32'bx;
            end
        endcase
endmodule